----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:51:55 03/11/2018 
-- Design Name: 
-- Module Name:    ALU_MUX - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity general_MUX_2_1 is
    Port ( X : in  STD_LOGIC_VECTOR (31 downto 0);
           Y : in  STD_LOGIC_VECTOR (31 downto 0);
			  Z : in  STD_LOGIC_VECTOR (31 downto 0);
			  W : in  STD_LOGIC_VECTOR (31 downto 0);
			  U : in  STD_LOGIC_VECTOR (31 downto 0);
           S : in  STD_LOGIC_VECTOR (2 downto 0);
           E : out  STD_LOGIC_VECTOR (31 downto 0));
end general_MUX_2_1;

architecture Behavioral of general_MUX_2_1 is

begin
process (X,Y,Z,W,U,S)
begin

if(S="000") then E<=X;
elsif(S="001") then E<=Y;
elsif(S="010") then E<=Z;
elsif(S="011") then E<=W;
elsif(S="100") then E<=U;
else E<=(others => '0');
end if;
end process;
	  
end Behavioral;

